PK   R�.U,�1�  �N    cirkitFile.json�]m��6��+�˳�5ե��[;��'��6�.�����1�س��I6�.e���Ԍ�{���f���#^�K�<�O?Ϛ�w�^��F/~��v�Y�n(�������~��g���b�Y����w����wo��^{E���p�E�	%5yYTU^XT�WP�yA��~��UY��n޼��7t�5�r�aq�Y��r��+o�pk�����Ha�#l|���X�ܼ�߬�z��"�*L�*��˰��2-�:�ˈB��a�gsWݠ�[�q�UQ�%-���˘�$��8-�ce<6m�6$�a��J��
˟��'����6>�;<��`���G����3���C,!�?i|�����������Y�PXzaru�^��K�<���(��9��K��n�M��6��gh|���_������X���6>���/q�'X�,��a�����S,)�?i|�������L����˟4>��G��x�.���7Xp�H�	"w�T1`��@ B+@`	���E �@�	"�C�.�+A����C$p���L�X"�"$��!8D�2�|a �,�q���!r��E�4�i�!8D��]&�j��X��H�	"w�\�!�bC`�F"�C$p��erن����q���!�%�nX�Q`�F"�C$p��er�F���n�!8D��]8��>��>�8>��n�\�Q`�F��q���!r�ɵ�nX��H�	"w�\�Q`�F��q���!r�ɵ�nX��H�	"w�\�Q`�F��q���!r�ɵ�nX��H�	"w�\�Q`�F��q��^�xd8)u]������בW$e�Q|�2�,��5���nz`��m����������U��ף����]'�{�9���r�0���i`��)q`�˱84Y��.�v������|�޲��GZ_�|�;����������-I��%>�/����kI=C�S����/L]kI?��0u�e��'�0�����5x�o�s�n�a/���u�/�u�=W(��Cɝ�Vc��.�y�ڪ���}��H)/K3e�ʼ<�K/)���
3�?����w��߹���{~�Pv�~����?��"�5{����q�(7�M#w�}�?��#�w�Q۝�u���y��t��1���� �2N.�fc��|��a�P�L��ÁaZ�8�|�G2
ڶꀣ�P�\����m�z�Q�L�(N.ߜ�Q�L����?�@��=Ea(����:���w��#'Smw`��Q�\�����m{{�Q�L'(N.���Q�L���]@�@�S'�o��@�AA�~!pT ���˷�pT Ӡ�mg8*R9��d�)��t�I�vX����Fc<,�o�Z6�\6�^F0������"��if���7���,'<,�o�r6I�#�0�����"���g���L�R�*xX$�0m���* �aB��C��E���&��a��&�Y�%xX$�0Em���- �a���m��E���&��a��&�Y.(xX$�0um��&0��*0}��K��"�����I�v�ŀ���k��
�7L_�$n���o܁��N�Mt$w&m�Ci��k
��Yn-xX$�0}m��f5 �a���낇E���&��ak���Y0xX$�0}m��8 �a�����E���&��a����Y�2xX$�0}m���: �a���?��E���&��a����YN5xX$�0}m��F=.��~= ��b�{ �c�5��g�M�}?����P�eN��u�p� Jǜ8�x�u���do�q��<�����&���p���A��Y��"_If=Lw��#�y0�,�PF�� `0Yܵ�aჀ���&������ �^�}{��-�K둾F:.���8ϯj���<�Q_���Q�z�<�/}MkL[.��;�}�B'Yw�����X¬�î�W�m��R���#9P�Y� �簄A��[�@8�^G�Q�L��vX Q�L+'֋h4*�iP�K4*�� ŉ�
�
d���
d:Dqb�|F���A���P�X��Ѩ@�AA;,aШ@�c'�g4*�iP�K4*��ŉ���
d���
d:Eqb�dF���A���P�X��Ѩ@�AA;,aШH�&���(pX�x��&��e	��'�M��M$��Բ��i�2�	f�5
�7L3�$n�%�o�lf[��a�|Ô�I�vY�`���g�5
�7L?�$n�%�o��f[��a�|�T�I�vY�`��	i�5
�7LK�$n�%�o��f[��a�|��I�vY�`���j�5
�7LW�$n�%�o��f[��a�|�ԵI�vY�`Ϋ��5��<���&��e	������(pX$�0}m��]�0�q�&:�6ё4ܙ���M��)��f[��a�|���I�vY�`���k�5
�7L_�$n�%�o��f[��a�|���I�vY�`���k�5
�7L_�$n�%�o��f[��a�|���I�vY�`���k�5
�7L_�$n�%�o��f[��a�|���I�vY�8`GX��Q:���0r��]�K9JǊp�%����5�F��1��X� `0��u\j�% ��]g�X� `09���l�%`��dq�z<� ���.	e�% ��]��1�0 L�,^��ޖ0rL[^P�-a�(/�ޖ0Ϣ�������QoK9ʋm�m	#G9m˗9���nQnV�f��>�n���ò����*/u�X��������A�%}�n�s��!Y�K��v�;KL&y�"�u�CV�Ĕܹ�%�� ��y������ L��a=ư@y��;��{���~�;�u��rM{o��\xҿ�����|�)V� �L+o�t�@8�� �~���k���+=m��O�n"���� G=� DHV�qŷ{X���~���ݸ;>,+���B�&�:W��ۿ�XHX%y�G Ľo���H��
I�N�
I%9	�F�BR��׭#�8<��V�8<���׭��8<��6�8<���׭�8<���8<��������3�BR�ÙBR#9	�>�BRcy�['/qx�!:�qxy�[�)qx�!:\qxSy�[�$qx�!:qx3y�[gqx�!:�	qxM  �؞|@@� Pw�Q�<�\���� �%Bԁ�:hY� ����p	�v�Q���\��'�� ���t� J�h<��%@�G����r)�=\�~@@� u�˿O�%@౽뀀.8J�7��K��c��1\�p�.�=)� ����b��=�(]�zR.���'�p	P}�Q���� ���Ĝ �>�(]^xR.����p	�}�Q�|�\"�����O� ������u�}l�6  �K�����O'�����l@@� ���{N�%@��}׀�.�8J����K��c{�1\tp�.�8)� ���Kb��>�(]~pR.����p	�}�Q��ޤ\t��������t����pp�Էv�#\�$��������ݒo�:�w|�w�$:�2¯MR�?c<�D ������qdX�1.l" i���x�� 2{`J<	ly��@���H3�^M ML{4�LM ML{�1�:M�L&��K��w|�ch�vL���z�m��o���C�/\�0S�����Aeo?��������NoK������j@8G�B�v�YVƫ��Ƭ��h�ݼ��6�5�`��~Ӌ1�I�O�2S�-hJ�)J�,��dJ�)N�<�
dj(SC�ئ�25���Lej(SC���L���W���sw��O�B�9�Ї��
Q�G��3O����t��y!U�I�%S��1�{2�zg�\�O���r�ǹ���1Rc;�� h�������H���	�f
�b�gO��X:��k���θe��B��H����G��2�n����/�K�})<\
�K��Rd_��|���W��I_/��f�Znw�TW�ERԩ�'�g83�I�yY��*�9/_ļ�]��y��W�X�zg7e��i�ze�'^Xq�UYz���ҾRil�����V�^�o�<ܛ��߁�x[
�bE�2gUW02ԧ���5ߙ'�������^7��n�����/�D���]�\������wsu>�=_=�߾3D����^rg������O�[Ɲ�Ԧ_��V7�,��b��>k�����f7;n)s�>_?�y�{h�awN���d�h	7�~�]��7�_�h����4��M��W\�WU�~�%Q�{	O/<8U��,�O�(	C3"x����N���|�i�LW�o̬M�rٔ+} ��J��h�(z7綪�0;�	/�I�@��|�|��|�]�>U��Ar�y<^�Tǅ��Fz^#�/d���
��F%s/ή�>IL�0�W..{�].I����X��O;/��ZAw���V�]ˢ�Y,��^Ŭ$q�s�]�N!w9;����s����Q�];6[�~�=T��/���-]ӵyL9fۋ�&�k�~F�y&��av�f����Fg3ON���X�?�CO�Q��❟zuT�~q9����\�<��׻�5�z�y�ڡgr*P������Qtm�Yz��)#x�LU�"��0�T��.�N)�_��Z�G1�{4��ix��qh��OG�Ҩ��C�Q�zVҏ�p����O������$�SG^�}��!?<���C/����a��A����y-ST^�ו��狺�������΃��9��Yx��!E�op0}Z���'H�謁n���W�����@�	��99YE�yz�IOӃ/&UP�r���#���Hi/����_�Vz��Kz�����t�G�,h'�����y�T��LGA2�7�J7��o[:��n�ζ��]y�v6;[V�'a�d��x�R�$�K&TVu�+}my��~�a�w�~�j_�']�7*5ߜ7;Q�e:$/2JҼt�u��O�Q�gQD���X+�W�G*��R�I��ޫ����r]�i�בǫ��#�{YY�W���2I�X�ܾZ�C��O�>��1�ۻ�:'�CUE��	x�*~`�)�5?�2��J����͛f���^�OP���S͹����y��4Kx�T�wy���f�O[��2�P�\ϲ:�¼��"�^��*�Kʋ�q���}����gFv0��������b�"��O�����W^o��wU����p�˜�t*��˕vd�5W:�(ޜT��8!t͏���2���Uy��.˴+�҂�6�� e
t�����-iUiTց+��(R��rO+��c�uyI��DU�Ұ;��¯��*��G���ν8�B�%�:γ�3����v��fY]m�����r������շ�^��>m���+S��N7z~��\5�O)7\���e�W��l�8������{��t��t
�o��z���S�|����~��?#����9�qx��L�_��V���tJ����O�O�t�5/+xGt�XJ�B�"�<^��Џ��Kx�� �$�u�	z�X���x,e�q�~���.��|��q+��|�g�y,q�ꗫ�n�����s��4g�X)�x���O=����m�K�g�>��|V�����B��e������ӽ�Jܚ"/���<��[�_:iԱ1�e��S�?�|���}^�G��c���г�F��n���I��鳰�f��y��D}�xl��"Z'�I�ny]���G���]Yރ+^&*��b�)��^���#�S?>�-�Q��P^d�W�F��bx1�9oD�X������~���Ҡ4��Ɂv0�6��3/;�%��y�9~�aY��L��x��nw:���n���~<���ۼ���;]}��8�n�n�闥��/�ߍ1��g�@�dj������Ou��jx�����o����u�,T��-T���4���u��%OM������ۙ��_�?�3��|z����Q�0D/΅S`ޖ��7۱��f>���ϱ�:���,�bg�Vd\���R����<}�9!S1¥bN���"�d��$P�N2Rg�ث�J���w�K�LE���W�T$\*R�E���y�d<ӛ;�lH���8ό^�<���y�3��5w%c{�_2�;��+��韋��#�n`*����9�l[�D&s|*�+f���q���;k�(^�c�ax�%<����(u|t,u���Q�k dA��u�A#�xq�zl��}(<��w+�bԚ�Tr�)A�N΋b�wn�(f���R�*uxx>ӟ�3t���%T��hS&T�7�4uhB��XWB]�2w�����[*�)�)
Cp��ۗ�;'8]�DG�Re@S�=봰c�yi�?w=���L��$�w�s�$�-�h����|�v%�E��=�����[�c�0b�r����!��f���w�9{��/����|����߼����K�7�̾�?PK
   R�.U,�1�  �N                  cirkitFile.jsonPK      =       