PK   ��9U�D^��!  y�    cirkitFile.json�]��6�}�F��^��(�K<l���H���(胊iW�TW��~�}�}��T��U�TE�=�����t������눺�c����y�Z���v}�X-g/(�����Շ|���rv�X�7��������������k�W��ՙE����#ʊ4���e
[FENJ�*�����ً�o/-ܬ>�u�����7��|����*�"�-��sc�a���X�z�Z��fnbk�eT�<�tV�Q�(�\ʈX�J9h��sbǊ��'l�������\�\b�'���C)U���Q��$҉5�1��D^R�%*I����e_ݴp=J���Uױ���\TQM�*-�un�k|���J�fsŎ���Fai��GX|���0���?��a�����������#,>�����	6~	6~���;��;�?s�6��k���id	S6kR,	S,	�������ܰ�`�g����#,>�����6~6~\|��GX|bN|݋����/6DC$0D�d 	�a�E,������:�,+Y���	��]��u%KV��	��]���%�K֗�	��]��5&�LV��	��]��&KM֚�	��]��k5k�	��]��+6�l�	��]��e�t��Q+��}���Q� Wb�M������ك���+F�I�bĆH`��蚌�I�b$��"�!�k���AqN�I���q�t)E�k������)��z.s���sS�S|�	��]���&	V�$XmbC$0DCtM�Yg� ��d&8�;B�/��p� ��_,|I��ņH`��蚌/|I��%��"�!�k���H˸�'X4�`�L�E3,DC�B��Ꞣ�r�M*���n!�i!�=	2��@�xA�]��^��wA�p�;��������y8�}�����]Ee�\ƫ����)��e��o4Mq�4�`��]��ޝ�GV��#�w{�X:s��?x����g������-���L�y�[��gҏ���*�Yq����bl}�PΤ�'ꍭϤ����Ϥ�����3� �E��{��s{�d�f?�&��<�
��4O�,�����,9��
�μ�p��>���$F��uR�����QF���d�����T}{P�a�AՇ����IRۨ2��")��d�eW�Vu&��AՏ`�
�,���kS���8y�m���">��!Շ�4]�=p�cl�(-�n=��4(���,x�����a��Yv���qs�~�{����Y+�8���]<�DGY,(*�XW:NM��u���Ý(0U�b�a�f,]���Ud&�K�~_�c{�&�T��^��y�f_����+���Sp����g��dT���Tp��Ә��11�J�[F�OA�
�.801�>�[F�]�pc2h?y&�
��%�U`�A���Rp��HkTL�'��V����3Q��#�b�=]�
�4���
n���	$�U`����,?�&�}��k���I#�U`�A��Rp��>mP1�'�[F�O6�
�t��I���*0� �~Z*�U`�	&�y���f��	L'�wO+P�qR�DZ�DbN-�H.�F/#�`�%�E���')�,2�0��K#�7��7L9�wO-P�a♗p
oo�~6	�|[�x�$4/5�,2�0m�=��@�	i^+�Yd�A�{�w��"��ӼtWx��x��Ip�d��&�y���f���j�����7LZ�Y;��k�Y�S���I�7�<��׼�Wx��#+0}m�=Y�@��k^�,�Yd�a��$�{��ә�Ze��Lt"m�#i0}m�=��@��k^�,�Yd�a��$�{��Q+/��,2�0}�7�,2�0}�ˀ�7��7L_�wO0P�a���+oo��6	�Ta�x�:S���*gf}�K��7L_�wOb0P�a���4O���p�$�E�;�f}��9���$L_���6;��)� V���	� VvY��q��u|&�>n�O�@40{�O��2���H��0�a��q�3�f!�l>�ȡ�0�����3k!̴,.�)��3�aX<���9a��!	�tZ3�#�ȱ�'���+�o7wF�+��}�š� V0���P�i��[	͎�r�]Bse��l���Y +��%0���I_B�j�Щy24O��ښ��:��MW՗Mb|ީ㻃ДQ�c�9ꄕ�R'&:��DN�c����cj��M����JK{�Y��<9�;܁���z���Z	�^Oj%�U�����w�mi��Jh��HKTL�h��H�@��VB[FZ�b��@[F�'��*0���*0� �=���V���Q1�o��#ݓZ	m����*0� �=���V��NQ1�l��#ݓZ	mi���wXmi��Jh��Hg��x�4�V����I����TN`"��bn)��t�Ip��V��'�M��M$��Բ��i�2�	f~�!�Yd�a��$��R+a����Cp��xÔ�Ip��V��&��)��f���g���K���7LB�S��"�S�&�ݗZ	o�����E���M��/�&�09�O17��7LQ�w_j%L�a���bno��6	��J�xä5?��,2�0um�}��0�U`���bnyd��M��/�&�0}�O17��7L_�w_j%L�q�&:�6ё4ܙ���M��I�����E���M��/�&�0}�O17��7L_�w_j%L�a���bno��6	��J�x��5?��,2�0}m�}��0��k~�!�Yd�a��$��R+a����Cp��x���Ip��V�����)��f���k���K��c���J|+�����VvYg�V�[X��Z�oe`�:#���@O;'����Cǥ�I�0�!�Й�sR+�`8<����J�Q��!����J 3I(�V���xhqNj%�����$��S+�`|9١�S+��Z�o�d��V�[9�.����VN�Khj%�����V�[��r�/����VNNK����Z	N�ķr2F����VN��Z�oeߗ��������j=_T��^��r�a����뼴�|���֕]�^�~�|8�Z����>�-)n�W:����tG���27�ľ�� :#x�m�k�y��eG�UP���
�8_��v�K��ҬbY7��`=�M��g����L�:�o���+�R�������U���{(���y�����n/�56+\UYW��*�ra\��β$)#�6])g�>��+Cn+]�(�����"�
aD��B��NY�#k���Ǭ��47BNC#e�p�O7�Ka+���3�`��{Q��[�&y\G����2��w�Yw�YН)c�z`p	�o� �Hi�{_0���l;� ��9����E<	�sn~Ns��fu�u-"�#��)��$5Ee�DAJ�����m���k��HW���*-�*���*-�H�̆����̛�*�&)\���!�BF���(O�I)��%3������Ѳ&m��L�te&ʲ8�
#H�"�I'�z�Ȁ+֝0�yp6�3|A(�փ��N����2�.R|*+�s���NL&Ar�ҙ�8��9��a��ѵy?&BΜl�a�������µ}���V�|Y�=7|��t����}އ�/�
H����R�W�'��W��{���}�����nP[eL���������C|?������'�O�{�x��|���蹝�L���O�(��Jg�{CT���E�'�3��������O*`�{�����|j:�{wzB���|���<6~�c��nFN���p����a�<�~��>����>�3���f�e&�1�l1^���B��O����q/����>������<�;��'r��Oq0�� �|.��1]��3:c׽O�>'+Or���\�"� }���$܁�$�c��&���@�9B�O����>�pN��K ��<�9�����'Ay�'�5�'Zi"|��N��i�3�҇���oL�C�a�cs�S���w��*��	�%�'x1!��ڳ��0B�?gT?g��H���|��%X�@,�A;�O�e�����@���	��"�����"��D��4%1G��uA�:�_R��?ɢ���$�B��E�ѧ�O�(�pp�)"|����^������v�o����ϫ���`�Y�������/fs�����F漡����5ҋ�8�C��M`���+�$�l��H`�����V��Њ������:sD`�F�����V�=HP�	����ؙ��}\gE6DC$0�m&|f�{�L�كD���	Q��)c���!T�=Ho��i��S!��{�vvL�����Ab̆H`��(گ�1[���)�$�l��H`����"�ս���A�ȆH`��(�_��������>JB�$4J���(���\�AH>p�-�@�!��Ch݇���(	�Rl?��mz��Ch�����(	�Rl�l�mz��Chч���(	�Rl?/�mz��Ch量��(	�Rl���mz��Ch����(	�Rl?��mz��Ch�����(	�Rl�v�mz��Ch�����(	��y���� �Q���
��	z�3f����@��# UH�U!�V��(	���(]�T!�V�$Z�$4JB�lӀx�%b	??��(	��5@$�h�H�E">JB�$4�6��M%3��2�}L��hi��$��DKH|��FIh��� �DKH-!�Q%�Q��ʼ��0�(I��$�%�Q���M�i-��>&� ��4�	m���)�	�y�^�I0Л�6 �	���f�
36?����Y��Ҍ�@�qR�΋{��#�y˅���9id}o�Y��?c�Ŧ'���!������5�m �����6� ���On�阾z=� {���W�����َ5�%��h����&<>O������Su��T�$��4*����<��LRdcH7+�,9���Ͻ��nT�H/IL�]R��I��J"#D��
����K{P�#����T����6IjUF4�1�"�HfQ]qUkUgB�T�����͒���8%��D�i[�8�����H�#�J�s���ɋC'��d[��2�5&0���3��	}t���'�rre��2N"��8�E��,�Y�+�&UG�T��s��Q1:wZ()��.0Q���/g�fU�}�ٿmү��f��gM�id��M3S7��f�m�7�6-ڐ��eԔ��(5e�)LM�6Y��A��G65dk��!��וeSC65�o8��i?p��n�}�,�E���b� �[1d�}���)`�<��G�C�����;����Bm��RE�&��FE�)�<Չ��(�
�u�\��3�z�%��n~ηf:��M���:�{'8ޡ?�yG�}���<�\џ��<T>çq<�b�G���t=��^�$ߞ��'�x�����x��"��]�񎙦�s&e����P���#�����y�W9�U�����_煽nj5ۨo�梹[��]�%�]"���]��%����K��R�]�{7�Ǐlw-�/��%�_Jv��R����~�$�"�W�vߑ_;>re��W����!���8���*�n^�n�D���ZW�*�-扚����;��Q�k[o�-�(��}�X_��?���7D��tPN�GӤm+=���W:��so;(��4s�_��w7Mj����޶��/�&ww���ի��Ʈ7��!��,����b�Y/��ȸ��7?7W/g���w�O_��k�v�\8�g��n߭>|�|���^����uo�������[��-ֶ���8�[���]�����]s`�؞'ۤ� O�+n�\l+��]�F\&���]c6�}�*�=nU�ͺ%�c�ڍ칐��r�I�T�f�p[�M�,�u�6ꗳ�zᢕo}�9�.�����u"��^rνN���g�IT 9TCՈ�j$C5���]��1��/�t����h�y0��.���2V�)��~o�L�����@y3P>(O4P��P=TÏ��񢸻�k�J~�v�`�.���]����������,6?l���'������+�&.�8���#77$��~��׿|}��uұ���.�61]�x�ܴFb�ǽ�$i���(SF�
+�(Qn�W�*Mk�����q�![�2�g���w))�j�O�-��ʤ� �+'���+�^P:��|f�iJ�Ӷ�2�#�v�#�O5��H�"�[[����J�Ed��vL�D�jA�p�Lg0j�pu�JN���v�z��n�J�����Kw���7=�����Ŷ��Q���=b��#���#��:lh�|[{Q}�/nxq����.k�Pr�G���qum�]�������ѧ�R�.�j"x��՝�b������?�O������O�b���^����}a���_�����ݲ{^8���$����C0�.�7�w�T�n�'n됫Hh�F�ۡE�T�uZ�_�v���!�N���6��Y|��4�W�3�������:��A�����a��?�J_�O�>�·Mi�	H�8�a����d䦽]O:X��D:ϋ:��Gq��Ȗq�2)ꢎ�R��
zv�m����w~�Eʭ��K�ۢYdE:K�t��v+Ou)U;ݹ��L[�5��L��,��n{�];�dȢnF�������l�\3�6�;fCv��I�x�� }��M�_}����|	_	F�1�6�0�Ζ.����wr��q�M�e�HEey]E������G�K���U�j�=O���Q��M��AJ�����Q�I��&ΗU^����o��]S��≤��u�l��P�Qf�b'��Z\�Uae�3��nS��n3�R�6us�ǣ��!<��#�XA�p��6R���G:�/�Y�;o�D��o�O_���_^^���lV�py�Դw��_=�e�7��4'A�������7/�%�W���ͻW�n+9o�������nY�\]�����L��#�/���q��տ���C�}7�/�p:j�y�5����=���9�u�Zn~X���Z}���8im�Ҟk/Ww�;�/�����]݈�*QnN�I�(���@n�L�H-�e�r]}�;���D2�U�E:Ү�F	չ�.�D��۝��=��Γ�n�7�)q�ڽ�\��ᜫvF��a	J���G(K)r7PW����@�!��Q����2�m��{/��v����zu]���oڦ3{�fv��ݔ���.��U�����JEi��a����t,���eR�㶼��ƍ
v�_����l�
��͓<��p���(��"�2JM^+�j�6�߫��By����f�/���,"i�̵�[l��z�,o�6{��ʘ2w�Ґ�tlE���[m��8/ӴL���7��mc�o�M��S���w��j�ZVq�vM!��\�j9-3�z�LӃ�x��׫�w7v�g��\��v�o$D.��:O"���E�67����zuk��ɵ"d��eu�p{Ѭrk	Q�\�n3���_�qe��k��7�Q��y ��?�ek�-���{Z�_y�Zo�������]�xI�Z��zqm{�t�*�3*֢�u�ak�����BFY��TIm��1�T�d��q!���L�����0YRPY�>F�8�����J�Q]���E����Q�oz�Q�uU�-{�zM���܂��ݶ�r�4�$ώ3����f��jQ]��������o�,/.���w����D��rє�xg���b��X�-/Vn�x�J��>n�i]�V�v��e�������V׿��z������#/���-��9��;J�bGOKO�Dͱ�f=�UwVn��EJ쌸��R��]Ln䊩=��aQm�5��|��;���]ҏ��V���~sn=/��꫇���v�������w7'���M���h}���Mն���v���g��2{Y��bnm��? }u��:��7��[M�w�qG�7��,�w������������́���xnh��M�˾Rio)���4��Rt��ۏn�t�<$��51�`�d[ڟ���$ؽ�c	���uJ%��Pr|���C�K�,`;�=�df�(��ot{WD��#�!���q~$庡��i"��R���44Ov��h�'�I��#i�9M�N���(�U�&�<B��/�Lp9W�~��cL��As�mt�X�ѠyΤr4R �	i��i��E���R:�/�3�J�R��n�^.q����щN��,�P���yl<x�m��6��J*���ل�,�eG�}քӦ�kf|!���;+�XH�6�P �Gm����.�����_�K�>w��<,q��c��P:>���#����ƾ	:G)U#|���g.�=.> �ТC�1�zHv(L�:\�K��dX.��#�^SO�N�#�˴�si�}{&-;�j�{H7����<�X�dg�+I��H����c��S�+g���;{R?�=� ����=���y=x�3�ձd>ܸJ�?2eg��p�<���SR���uE�w�-%�R��a���g��G�
v������e�DC�*zh�P^�1�A!l]��b�A@���Y���	Z�vJl�TsL K)�G7v�b�G�;��a����+��1*,�ɔ�:1���*�QC�HG�yThh5Ҝ�Y\_W�-���"�n�W��s��������/���V�����!��o?�>�PK
   ��9U�D^��!  y�                  cirkitFile.jsonPK      =   �!    