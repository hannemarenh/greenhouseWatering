PK   �9U���  �@    cirkitFile.json��n�F��_%P0w��*���dv��LI�����naԒW���6���e������2�hS�~�d��@�m�uX��WE�:�4ٕ�֛�b��g�ֻ�j��\�d:y_����tr����ٻ]y�~r���~�����.��ִ�euU,cU�\� �t�J-����U�u��pN�o���o?ֻ`W�ֽ����r�:�n�'wS�gC�a����Lg��.�jZ�!�'�Δ�C�����O�O���/��g�m��p��ԛ�l�Q��"(�j�y��\A���E��"�G3]'�f�׬�Z,�O���Y$���/b���S,?��g�x�cV���O�O���/�%���Kȋ���QH�Xygt08��R��Mم e���S,?��g��",N���>c���b���/����Y�rV?)?��S,�pV��`�+X����O���:4�0`JLQ�L��C�F�DV�E�f��:.V���LQ�͐�}%K
v��LQ�͐��%�K
���LQ�͐I���;b�
��`�f����[<b�
��`�fȤV���U��1EST0E3dr�F����-1EST0E3dr�F�����1EST0�p��ލ��{7b�
��`�f��ލ��{7b�
��`�f��ލ�_��^����-�n4��hػST0ES4C&�n4��hػST0ES4C&�n4��hػST0ES4C&�n4��hػST0ES4C&�n4��hػST0ES�R�Q��{7b�
��`���ցx�c�	����b�W OdpWT6��2rG��s���j{)����y������ۖ��T��y[XAW�}6o_m\ؼ}���y{}��y{�]Z��ְ��ʥ�U�<�������ǔ�/��4�롤/�Rv0\�
k�1U/m/�e�H��������K�kٹa����oe��o�uD����G�ڏ�k?N�i��i�,uċ�"�U,�b��:�a�P��£wO�^ͻ�]Z�uZ$Q��Ԍ]��(�� ���$��*
���j�ͽW�nws�EZ��<P*3͋�
�EI��*_�a}�{������2��t,�eĪ\EnfN��j>_�:O��ޫys��M{���خ�;y���7oB�g"��k?c�Q���ɷa�F�I��GS��&��螛W���JC��TZ7@u�(�L���ZF��[FiMi2i7��Q:�4i?��QA�!�n��
*S����⨠�i7G�N�k��saT:�4qIè��)5��ώqTPi���h���Jg���0�e���/3J��23Jg�&c�vc,�sJ��3hT"�&]ਠ��I��1�
*�v31pT�9��"OPK�'�O6
oO��7g��䕍d�qn�Hv�8~���#O�K�yf���s@zc���a�Òzc��(�=�ޘy�]�ޘ6
oO��7�&y�?xXRo�E��'�3Ҝ����F��	��%O�K�9j���D�@zc�����Òzc��(�=�$�ޘ���w�ޘ�6
oO|	��
�9I<,��
母��t��kN&K��k���D�@zc����Òzs懶�R�8����5'g��%����Qx{bV �1�I$�aI�1mޞ@Ho�_s�KxXRo�_��'���ל�����F��	y����5'��%����Qx{�` �1�IN�aI�1mޞ�Ho�_s�N�w̝���,��k�4l�ޗG� (���0 J�]��q0�b�<��K�u��. Jǚxy�QuP�2����Ԁ���s@Ô����Z? ؅�S�]6������.�k@�Tq�߀\��b�[Cr^&���l!NޯVq�� ��˫�o���(}�] �Wǥo�����}P^��!0 �y_�"a���P�0���+ײ�8�4�z�G����牄�Q1��HD�q4�
*��D�Ш�Қ��yM��JC�=�04*�tDi�<��QA�!ҞHT:�4q>Ө��iO$�
*�P�8��iTPi��'�F�N)M��4*�4D�	C��Jg�&ΣfT"퉄�QA�sJ�!3�
*��D�Ш�����x�F��H{"ahT�9�L27�%��'��/�ћ��F��F2�8�l$�l�La����Òzc��(�}�0�ޘm�F�తޘs6
o_$�7f���(8,�7柍��	��Yhn4
Kꍹh���E�0zcF���Òzc^�(�}�0�ޘ��F�తޘ�6
o_$�7f���(8,�7櫍��	��Ykn4
Kꍹk���E�0�`����Ò��`��(�}�0�ޘ��F�తޘ�6
o_$�7�B�Ho���J�N�H/���i�_s�QpXRo�_��/�����h����F�틄a���57�%����Qx�"a�1͍F�aI�1m޾HFo�_s�QpXRo�_��/�����h����F�틄a���57�%����Qx�"a<�"a�(�ŀH9J�]րH9J��H9J��k@$��c���`���z]jH$ �p�;C"a ������V=�����!�0 S�]ʐH �����!�0 S�S�ѫU�;F�����	�;�E�ޑ0r�Wǥw$���q�	#Gyu\zG��Q���yj~��0[l���lU�6������]��ݯ�E]�V��vWջ��͍�֬��YtN�$`g���O����7�f�H���?n�c�=�tEe\_��pw������_�
Rn*�brczmv���iEE�/��>}���Ӊ���6]?���d�X����u�NHO>��A��"{22�<�6_B���].������
�C[dt�W3G�?>2����m ��(�E]�d rx��b���CQQ�S).<���ەBQ�\��'�P(j$u��IQQL�\��!*��Qw^����=���b�.�J&����h��Ɖ\�1��h��g��j#���(����3w*i����BQ���frX��<A���|ԝ�9<DE1EOb ���X�G�yא�CTS��rx�c vE|�  c ��җ�'Ւ�p�7���hH�-_f�h	?0K_6�TK��qs�@@FK���Y�r��Z��92Z&�җ�'�Rl��r�@@FK��Y���Z~��2Z��җ�'�R����@@FK��Y�r�Zf���2Z~�җa'��|��6��p}`��|:�;���f����{����e�I�|7wd�|��/WN�%����j  �%������h��q��@@FK���Y���Z����2Z��җ�&��}ܜ3���}`��7�����f���������e�I�|7�d�|��/M�%����c  �%���,}�jR-���k��~��H����\!w@@����$���j���}Ȁܴ��r@���;�)@h�����J����龝2$M�܏	AH�Py^�N$xҺt��!�g" �J)-L׳�n&��{K4$�L���-�������k&:��P����$��a��N.�h�;�L����s�$�_��;�L������$���<�<�[U6�� �mC�i4����$�@�<�)m�+�I05��L	b#XT���S�]��Wٝ��[�ݛ
e(�B����-�m�mm[h�B�M�J��fjߙn��n�M�>��m�G����A����m�Uhf6�ֲ�&��M:+�����t|�{���cs���C�5����ϓ|��.��O�y�����.����]w�N�Q��Sݝ/�&�nҧM���6E���)v7%�M�=1�����V��v�^�v|#��t�Z�55��0��Ea�<YF:�Th��M��~�=���,�������d>��ë�8��sy}�<�:ۭ޽?�R����Rb�+������n{_���9�~���lY�1�v��;3����n�N~-����������Y��O�O��ۏ?l�fp'��r����}��e�_�����v�>�vu5�>"F���aY.;��݁���zr�kzb�b���ښq�Iԕ>�x�&�Ub���{�Ȝ�y�Q�%Idq��P�͜��'Y�ű-{s�r(7�c�^�,��v�2j�ǾL��G��n��O��D����4û�M��?O;��:�/:�WaG��ZD]-Ү��J.Z;ŧZ���E�jq�<��.Q��9}>�t~ڐ���O�����y�np�<��?��?�ؿ��_��NG��W�ӆF��Ϯ>��q�9mp�9mp����5������C���R���I���UhNҥ��?*���O���t_����a��f:ϯ�6���Fx�����c���-/��<[��-���������yPG*��4�TU�^�z���X�t��O�t��f{6��9�}�r�s/TWy��*�ڮ��<��49?��*�4� �WZ��RjK�U�:ȣ|�uXy΃4J��
�,[F�R�uܣԜ��Ti���_IZ��J����k��Tq��q܏�~u�3ѫ���g;=I�lo�����n)n�l�۴^U?��w��Ef�\�$���1�b�~ޮ�]�G������OO{=u)��U��
�ol�+�|^��?�o����u�5������3G���a^��a��w�ڿؿ��g�|�Is������|bxjJ��-:��^���$�ei*=�� I�$�U���l�/��Y��<�q�Mxun���cm��׻_>�����?Z�ͩ����W��z��?���Su�x%ѫL����qx���R;�s��1��*���:��#&Wf͏�]������ˎ��[������}]}��2x����Y���F�۪�t;i������ɷo�ئ��魹(w�����U�Ib�6x���I��zW~������y`>���������v�9�-��O�������|k7��\����7�o{�����T�-�v��o/�������)�� ~���|%�^|O�/�^�.~{���u�5,~���?7O�l�_V{X_/��^�	�C���U�x��_*�#��+QI��
�xQ*��4XP�x��*�����R��{u��5�.ޫoA�8=]��=7��۽V]��
��|ݽ���g:���i���nv
Ԡ�ܓ�i�h���}K�
S/���^�;uv�{�屢X��Z1uw���J'�N�M���ܰ�/g�c}ٛ��z�����ޭ�}��A3%�o~Y�W]���<����?���������PK
   �9U���  �@                  cirkitFile.jsonPK      =   �    